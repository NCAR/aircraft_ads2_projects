THDR       h3.0     278     0                                           N312D      \  �     '\ADS     HDR        $                       SDI        p         2  QCW     A      :�M   BP	7���o                                                    SDI        p         2   TTRF    A      :�M   �~(��L0:ѷ                                                SDI        p         2  SPARE1  A      :�M       ��                                           �P       SDI        p         2   QCR     A      :�M   BN�����:��IR                                                SDI        p          2  TTB     A      :�M   �$b��8�	�'                                                SDI        p   "      2   VLA     A      :�M       ��                                                      SDI        p   $      2  ADIFR   A      :�M   =��2@�49ѷ                                                SDI        p   &      2   BDIFR   A      :�M   ��7�@��j;K)_                                                SDI        p   (      2  AVZI     D      ?�         ?�                                                      SDI        p   *      2  BPHDG    D      ?�         ?�                                                      SDI        p   ,      2  BROLL    D      ?�         ?�                                                      SDI        p   .      2  BPITCH   D      ?�         ?�                                                      SDI        p   0      2  NCNTS    D      ?�         ?�                                                      SDI        p  ,        FMRB    A      L:�M   �#�
B�O�=���                                                SDI        p  .         FMRR    A      L:�M   ��/BzL�<-�                                                SDI        p  0        FMT     A      L:�M   �>�RBD<[��                                                SDI        p  2         FMB     A      L:�M   >��uB��F����                                                SDI        p  4        TTFH    A      L:�M   �   ��                                                      SDI        p  6         FCN     A      L:�M   =m�h�A�                                                    SDI        p  8        PCN     A      L:�M   @E��  ��T�                                                SDI        p  :         XICN    A      L:�M       ��                                                      SDI        p  <        VDET    A      L:�M       ��                                                      SDI        p  >         VIT     A      L:�M   ����!J#                                                    SDI        p  @        VTH     A      L:�M   <#�
�!��                                                    SDI        p  B         VDT     A      L:�M   ==�|��q,                                                    SDI        p  D        LWC     A      L:�M       ��                                                      SDI        p  F         PLWC    A      L:�M       ��                                                      SDI        p  H        DPT     A      L:�M   ��u�Xy����                                                SDI        p  J         DPB     A      L:�M   ={���8:�-�                                                SDI        p  L        	CO      A      L:�M       �L��                                                    SDI        p  N         	CMODE   A      L:�M       ��                                                      SDI        p  P        
PSW     A      L:�M   Dj��Y-;ě�                                                SDI        p  R         
VDTER   A      L:�M       ����                                                    SDI        p  T        TEO3    A      L:�M       ��                                                      SDI        p  V         HGM     A      L:�M   C�s3��                                                    SDI        p  X        FMRT    A      L:�M   ?b�\B�G�=�v�                                                SDI        p  Z         FMRL    A      L:�M   >��B��;��>�                                                SDI        p  \        DTT     A      L:�M   �C(�@���>+�V                                                SDI        p  ^         STT     A      L:�M   �F�@���>,�                                                SDI        p  `        DTB     A      L:�M   �N�@���>1&�                                                SDI        p  b         STB     A      L:�M   �Ly>@��>/�W                                                SDI        p  d        TWET    A      L:�M       ��                                                      SDI        p  f         TDRY    A      L:�M       ��                                                      SDI        p  h        RICE    A      L:�M       ��                                                      SDI        p  j         IRT     A      L:�M   D�h��sLͿ�1�                                                SDI        p  l        IRB     A      L:�M   D��RÆ�����                                                SDI        p  n         SPARE2  A      L:�M   D�vf��33��PH                                                SDI        p  p        BCROLL   D      L?�         ?�                                                      SDI        p  r        EPSFD2   D      L?�         ?�                                                      SDI        p  t        EPSFD    D      L?�         ?�                                                      SDI        p  v        FETORQ   D      L?�     D��>2�x5��                                                SDI        p  �        HTWCH1   D      ?�         ?�                                                      SDI        p  �        HSDWP1   D      ?�         ?�                                                      SDI        p  �        HTWDB1   D      ?�         ?�                                                      SDI        p  �        HSDWC1   D      ?�         ?�                                                      SDI        p  �         HTWDA1   D      ?�         ?�                                                      SDI        p  �        NTET     D      ?�     �B�;�l�Ψ�                                                SDI        p  �        NTEP     D      ?�     B�=�CB4�a�                                                SDI        p  �        VUWY2    D      ?�         ?�                                                      SDI        p  �        VUWY     D      ?�         ?�                                                      HSKP       p  �        �V10     A       :�M       ?�                                                      HSKP       p  �        �V10R    A       :�M       ?�                                                      HSKP       p  �         �TADS    A       ;�`W       ?�                                                      HSKP       p  �        �TV10    A       ;�`W       ?�                                                      HSKP       p  �        �FLOADS  A       ;�`W       ?�                                                      HSKP       p  �        @�FZV     A       :�M       ?�                                                      HSKP       p  �        ��FZVR    A       :�M       ?�                                                      HSKP       p  �        �VDREF   A       :�M       ?�                                                      HSKP       p  �        �XV10    A       :�M       ?�                                                      HSKP       p  �        @�XFZV    A       :�M       ?�                                                      HSKP       p  �        $�VP15D   A       ;ps�       ?�                                                      HSKP       p  �        4�V28     A       ;�z�       ?�                                                      HSKP       p  �        �VP15A   A       ;ps�       ?�                                                      HSKP       p  �        �VM15A   A       ;ps�       ?�                                                      HSKP       p  �        (�TEMP1   A       ;�`W       ?�                                                      HSKP       p  �        8�TEMP2   A       ;�`W       ?�                                                      HSKP       p  �        (�TMP1    A       :�M       ?�                                                      HSKP       p  �         �TA2D    D       ?�         ?�                                                      HSKP       p  �        �TS2D    D       ?�         ?�                                                      HSKP       p  �        �TLSI    D       ?�         ?�                                                      DIGOUT     p  �         tDOUT1   D       ?�         ?�                                                      DIGOUT     p  �         uDOUT2   D       ?�         ?�                                                      SDI        p  �          DUMMY   D                                                                          PMS1D      8  �   �      h   `FSSP    IBR             PMS2D      4    �2D-P    IBL     2DP10           PMS2D      4    2D-C    OBL     2DC18           PMS1V2    <  �  X   
  
   A           FSSP    FSTB    FRST    FACT    FSTT    FTMP    FANV    FSIG    FREF    DUMMY   DUMMY   DUMMY   DUMMY       ?�          ?�          6v��        ?�      A�p����ɴ�F:ѷ8��    :�҉8���    <��{:S��        ?�          ?�          ?�          ?�      OBR     FSSP122         PMS2D      4  �   2D-G    OTH     2DGA218         INS        (     �   �  A  A        GPS        $  �   D                LRNC       $  �   �                